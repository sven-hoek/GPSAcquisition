`ifndef INCLUDE_ULTRASYNTH
`define INCLUDE_ULTRASYNTH
 
  `define RUN_COUNTER_WIDTH 10
  
`endif // INCLUDE_ULTRASYNTH
